6#3